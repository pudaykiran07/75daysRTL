module mux16_1_tb();
reg [0:15] in; 
reg [0:3] sel; 
wire out;

mux16_1 dut(in,sel,out);

initial
begin
#20 in=16'b1000000000000000; sel=4'b1111; 
#20 in=16'b0100000000000000; sel=4'b0001; 
#20 in=16'b0010000000000000; sel=4'b0010;
#20 in=16'b0001000000000000; sel=4'b0011;
#20 in=16'b0000100000000000; sel=4'b0100; 
#20 in=16'b0000010000000000; sel=4'b0101; 
#20 in=16'b0000001000000000; sel=4'b0110;
#20 in=16'b0000000100000000; sel=4'b0111;
#20 in=16'b0000000010000000; sel=4'b1000;
#20 in=16'b0000000001000000; sel=4'b1001;
#20 in=16'b0000000000100000; sel=4'b1010; 
#20 in=16'b0000000000010000; sel=4'b1011;
#20 in=16'b0000000000001000; sel=4'b1100; 
#20 in=16'b0000000000000100; sel=4'b1101; 
#20 in=16'b0000000000000010; sel=4'b1110; 
#20 in=16'b0000000000000001; sel=4'b1111;
end 
endmodule
